`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/29/2022 04:32:34 PM
// Design Name: 
// Module Name: ROM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define ADDR_WIDTH 5
module ROM(  
input [`ADDR_WIDTH-1:0] i_addr_in,
output [23:0] o_data
 );
 
 
 
 
 reg [23:0] mem[0:31];
 assign  o_data = mem[i_addr_in] ;
     
     
 initial
    begin
      mem[0] = 24'b00111100_01010101_10101010 ;
      mem[1] = 24'b00100100_01000101_10101011 ;
      mem[2] = 24'b00111100_10000101_10000010 ;
      mem[3] = 24'b00000100_00010101_00001010 ;
      mem[4] = 24'b00000110_01010101_00101011 ;
      mem[5] = 24'b11111101_00010101_00101010 ;
      mem[6] = 24'b10101000_11110000_10101011 ;
      mem[7] = 24'b00111100_01010101_00111011 ;
      mem[8] = 24'b10111101_11011101_10101110 ;
      mem[9] = 24'b00111101_01010001_00101011;
      mem[10] = 24'b01101100_11010011_10101010 ;
      mem[11] = 24'b10010100_01010101_10101011 ;
      mem[12] = 24'b00111100_11010101_10101010 ;
      mem[13] = 24'b1000100_01010101_10000011 ;
      mem[14] = 24'b00100100_01010000_10101010 ;
      mem[15] = 24'b10111100_01010101_10001111 ;
      mem[16] = 24'b00001101_01011101_00101010 ;
      mem[17] = 24'b10110000_11010101_00111011 ;
      mem[18] = 24'b00110100_01010101_10111110 ;
      mem[19] = 24'b10101100_11011101_11111011 ;
      mem[20] = 24'b001101100_01011101_10101010 ;
      mem[21] = 24'b10110100_11010101_11101011 ;
      mem[22] = 24'b00001100_01110101_10111010 ;
      mem[23] = 24'b10110100_11011101_00101011 ;
      mem[24] = 24'b00101100_01110101_10111010 ;
      mem[25] = 24'b10101100_1010111_00111011 ;
      mem[26] = 24'b00110100_01011001_10101010 ;
      mem[27] = 24'b00111000_11110101_00111011 ;
      mem[28] = 24'b10101100_11011101_10101010 ;
      mem[29] = 24'b000011100_10010101_00111011 ;
      mem[30] = 24'b10111100_01011101_10111010 ;
      mem[31] = 24'b0011100_01000101_00111010 ;
    end  
     
     endmodule 
